library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity uart_rx is
    port (
        clk         : in  std_logic;
        rx_line     : in  std_logic;
        
        -- Output 32-bit Integer
        data_out_32 : out std_logic_vector(31 downto 0);
        
        -- Valid Pulse
        data_valid  : out std_logic
    );
end uart_rx;

architecture behavior of uart_rx is

    component uart_rx_byte is
        port (
            i_CLOCK         : in  std_logic;
            i_RX            : in  std_logic;
            o_DATA          : out std_logic_vector(7 downto 0);
            o_sig_CRRP_DATA : out std_logic;
            o_BUSY          : out std_logic
        );
    end component;

    signal s_rx_data    : std_logic_vector(7 downto 0);
    signal s_busy       : std_logic;
    signal s_busy_prev  : std_logic := '0';
    
    signal r_buffer_32  : std_logic_vector(31 downto 0) := (others => '0');
    signal r_byte_count : integer range 0 to 4 := 0;

begin

    inst_uart_byte: uart_rx_byte
        port map (
            i_CLOCK         => clk,
            i_RX            => rx_line,
            o_DATA          => s_rx_data,
            o_sig_CRRP_DATA => open,
            o_BUSY          => s_busy
        );

    process(clk)
    begin
        if rising_edge(clk) then
            
            data_valid <= '0';
            s_busy_prev <= s_busy;
            
            -- Detect Falling Edge of BUSY (Byte finished)
            if s_busy_prev = '1' and s_busy = '0' then
                
                -- Shift Left and Insert New Byte
                r_buffer_32 <= r_buffer_32(23 downto 0) & s_rx_data;
                
                if r_byte_count < 3 then
                    r_byte_count <= r_byte_count + 1;
                else
                    r_byte_count <= 0;
                    data_valid   <= '1';
                    -- Use assembled buffer + new byte for final output
                    data_out_32  <= r_buffer_32(23 downto 0) & s_rx_data;
                end if;
            end if;
            
        end if;
    end process;

end behavior;